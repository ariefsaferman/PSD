library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
 
entity full_adder is
  port (
	 i_carry : in std_logic;
    i_bit1  : in std_logic;
    i_bit2  : in std_logic;
    o_sum   : out std_logic;
    o_carry : out std_logic
    );
end full_adder;
 
 
architecture behaviour of full_adder is
 
  signal w_WIRE_1 : std_logic;
  signal w_WIRE_2 : std_logic;
  signal w_WIRE_3 : std_logic;
   
begin

	W_WIRE_1 <= i_bit1 xor i_bit2;
	W_WIRE_2 <= i_bit1 and i_bit2;
	W_WIRE_3 <= W_WIRE_1 and i_carry;
	o_sum <= W_WIRE_1 xor i_carry;
	o_carry <= W_WIRE_3 or W_WIRE_2;
  
end behaviour;